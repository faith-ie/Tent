module tent;
  initial 
    begin
      $display("    _____________________\n   /                   / \\        z\n  /                   /   \\      z\n /                   /     \\    z\n/                   /       \\  z\n___________________/---------\\\n");
      $finish ;
    end
endmodule
